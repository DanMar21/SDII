LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY INVERSOR IS
PORT(I: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		O: OUT STD_LOGIC_VECTOR(3 DOWNTO 0));
END INVERSOR;

ARCHITECTURE STRUCTURE OF INVERSOR IS
BEGIN
	O(3)<= NOT I(3);
	O(2)<= NOT I(2);
	O(1)<= NOT I(1);
	O(0)<= NOT I(0);
END STRUCTURE;
